module bkadder(CLK, RST_N, A, B, CIN, COUT, S);//16 brent kung adder
  //inputs
  input CLK, RST_N;
	input [15:0] A, B;
  input CIN;
  //outputs
  output reg [15:0] S;
  output reg COUT;
	//intermediate values
	reg [15:0] B_reg;
	reg [15:0] A_reg;
	reg CIN_reg;
	//start level
	reg [15:0] p;
	reg [15:0] g;
	//-------------------------------------------------------------------------------
	//level 1 outputs
	reg G15_14;
	reg G13_12;
	reg G11_10;
	reg G9_8;
	reg G7_6;
	reg G5_4;
	reg G3_2;
	reg G1_0;
	
	reg P15_14;
	reg P13_12;
	reg P11_10;
	reg P9_8;
	reg P7_6;
	reg P5_4;
	reg P3_2;
	reg P1_0;
	//-------------------------------------------------------------------------------
	//level 2 outputs
	reg G15_12;
	reg G11_8;
	reg G7_4;
	reg G3_0;
	
	reg P15_12;
	reg P11_8;
	reg P7_4;
	reg P3_0;
	//-------------------------------------------------------------------------------
	//level 3 outputs
	reg G15_8;
	reg G7_0;
	
	reg P15_8;
	reg P7_0;
	//-------------------------------------------------------------------------------
	//level 4 outputs
	reg G15_0;
	
	reg P15_0;
	//-------------------------------------------------------------------------------
	//level 5 outputs
	reg G11_0;
	
	reg P11_0;
	//-------------------------------------------------------------------------------
	//level 6 outputs
	reg G13_0;
	reg G9_0;
	reg G5_0;
	
	reg P13_0;
	reg P9_0;
	reg P5_0;
	//-------------------------------------------------------------------------------
	//level 7 outputs
	reg G14_0;
	reg G12_0;
	reg G10_0;
	reg G8_0;
	reg G6_0;
	reg G4_0;
	reg G2_0;
	
	reg P14_0;
	reg P12_0;
	reg P10_0;
	reg P8_0;
	reg P6_0;
	reg P4_0;
	reg P2_0;
	//-------------------------------------------------------------------------------
	//carry level
	reg [16:0] C;
	//-------------------------------------------------------------------------------
	//output level
	reg [15:0] S_int;
	//-------------------------------------------------------------------------------
  
  always @(A_reg or B_reg or CIN_reg) begin
	//starting level
	g = A_reg & B_reg;
	p = A_reg | B_reg;
	//-------------------------------------------------------------------------------
	//level 1
	//generates
	G15_14 = g[15] | (p[15] & g[14]);
	G13_12 = g[13] | (p[13] & g[12]);
	G11_10 = g[11] | (p[11] & g[10]);
	G9_8   = g[9]  | (p[9]  & g[8] );
	G7_6   = g[7]  | (p[7]  & g[6] );
	G5_4   = g[5]  | (p[5]  & g[4] );
	G3_2   = g[3]  | (p[3]  & g[2] );
	G1_0   = g[1]  | (p[1]  & g[0] );
	//propagates
	P15_14 = p[15] & p[14];
	P13_12 = p[13] & p[12];
	P11_10 = p[11] & p[10];
	P9_8   = p[9]  & p[8] ;
	P7_6   = p[7]  & p[6] ;
	P5_4   = p[5]  & p[4] ;
	P3_2   = p[3]  & p[2] ;
	P1_0   = p[1]  & p[0] ;
	//-------------------------------------------------------------------------------
	//level 2
	//generates
	G15_12 = G15_14 | (P15_14 & G13_12);
	G11_8  = G11_10 | (P11_10 & G9_8);
	G7_4   = G7_6   | (P7_6   & G5_4);
	G3_0   = G3_2   | (P3_2   & G1_0);
	//propagates
	P15_12 = P15_14 & P13_12;
	P11_8  = P11_10 & P9_8;
	P7_4   = P7_6   & P5_4;
	P3_0   = P3_2   & P1_0;
	//-------------------------------------------------------------------------------
	//level 3
	//generates
	G15_8 = G15_12 | (P15_12 & G11_8);
	G7_0  = G7_4   | (P7_4   & G3_0 );
	//propagates
	P15_8 = P15_12 & P11_8;
	P7_0  = P7_4   & P3_0;
	//-------------------------------------------------------------------------------
	//level 4
	//generates
	G15_0 = G15_8  | (P15_8 & G7_0);
	//propagates
	P15_0 = P15_8  & P7_0;
	//-------------------------------------------------------------------------------
	//level 5
	//generates
	G11_0 = G11_8  | (P11_8 & G7_0);
	//propagates
	P11_0 = P11_8  & P7_0;
	//-------------------------------------------------------------------------------
	//level 6
	//generates
	G13_0 = G13_12 | (P13_12 & G11_0);
	G9_0  = G9_8   | (P9_8   & G7_0);
	G5_0  = G5_4   | (P5_4   & G3_0);
	//propagates
	P13_0 = P13_12 & P11_0;
	P9_0  = P9_8   & P7_0;
	P5_0  = P5_4   & P3_0;
	//-------------------------------------------------------------------------------
	//level 7
	//generates
	G14_0 = g[14]  | (p[14]  & G13_0);
	G12_0 = g[12]  | (p[12]  & G11_0);
	G10_0 = g[10]  | (p[10]  & G9_0);
	G8_0  = g[8]   | (p[8]   & G7_0);
	G6_0  = g[6]   | (p[6]   & G5_0);
	G4_0  = g[4]   | (p[4]   & G3_0);
	G2_0  = g[2]   | (p[4]   & G1_0);
	
	P14_0 = p[14]  & P13_0;
	P12_0 = p[12]  & P11_0;
	P10_0 = p[10]  & P9_0;
	P8_0  = p[8]   & P7_0;
	P6_0  = p[6]   & P5_0;
	P4_0  = p[4]   & P3_0;
	P2_0  = p[2]   & P1_0;
	//-------------------------------------------------------------------------------
	//carry level
	C[0]  = CIN_reg;
	C[1]  = g[0]   | (p[0]   & CIN_reg);
	C[2]  = G1_0   | (P1_0   & CIN_reg);
	C[3]  = G2_0   | (P2_0   & CIN_reg);
	C[4]  = G3_0   | (P3_0   & CIN_reg);
	C[5]  = G4_0   | (P4_0   & CIN_reg);
	C[6]  = G5_0   | (P5_0   & CIN_reg);
	C[7]  = G6_0   | (P6_0   & CIN_reg);
	C[8]  = G7_0   | (P7_0   & CIN_reg);
	C[9]  = G8_0   | (P8_0   & CIN_reg);
	C[10] = G9_0   | (P9_0   & CIN_reg);
	C[11] = G10_0  | (P10_0  & CIN_reg);
	C[12] = G11_0  | (P11_0  & CIN_reg);
	C[13] = G12_0  | (P12_0  & CIN_reg);
	C[14] = G13_0  | (P13_0  & CIN_reg);
	C[15] = G14_0  | (P14_0  & CIN_reg);
	C[16] = G15_0  | (P15_0  & CIN_reg);
	//-------------------------------------------------------------------------------
    //output level
	S_int = (A_reg ^ B_reg) ^ C[15:0];
	S <= S_int;
	COUT <= C[16];
  end
 
	//Registering the data in and out on posedge of clk
	always @(posedge CLK or negedge RST_N)
	if (RST_N == 1'b0) //Active low reset because of the std cell library
	begin
		A_reg <= 16'b0;
		B_reg <= 16'b0;
		CIN_reg <= 1'b0;
		S <= 16'b0;
		COUT <= 1'b0;
	end
	else
	begin
		A_reg <= A;
		B_reg <= B;
		CIN_reg <= CIN;
		//S <= S_int;
		//COUT <= C[16];
	end
endmodule
