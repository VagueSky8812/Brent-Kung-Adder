module bkadder (CIN,
    CLK,
    COUT,
    RST_N,
    A,
    B,
    S);
 input CIN;
 input CLK;
 output COUT;
 input RST_N;
 input [15:0] A;
 input [15:0] B;
 output [15:0] S;

 wire \A_reg[0] ;
 wire \A_reg[10] ;
 wire \A_reg[11] ;
 wire \A_reg[12] ;
 wire \A_reg[13] ;
 wire \A_reg[14] ;
 wire \A_reg[15] ;
 wire \A_reg[1] ;
 wire \A_reg[2] ;
 wire \A_reg[3] ;
 wire \A_reg[4] ;
 wire \A_reg[5] ;
 wire \A_reg[6] ;
 wire \A_reg[7] ;
 wire \A_reg[8] ;
 wire \A_reg[9] ;
 wire \B_reg[0] ;
 wire \B_reg[10] ;
 wire \B_reg[11] ;
 wire \B_reg[12] ;
 wire \B_reg[13] ;
 wire \B_reg[14] ;
 wire \B_reg[15] ;
 wire \B_reg[1] ;
 wire \B_reg[2] ;
 wire \B_reg[3] ;
 wire \B_reg[4] ;
 wire \B_reg[5] ;
 wire \B_reg[6] ;
 wire \B_reg[7] ;
 wire \B_reg[8] ;
 wire \B_reg[9] ;
 wire CIN_reg;
 wire \C[16] ;
 wire \S_int[0] ;
 wire \S_int[10] ;
 wire \S_int[11] ;
 wire \S_int[12] ;
 wire \S_int[13] ;
 wire \S_int[14] ;
 wire \S_int[15] ;
 wire \S_int[1] ;
 wire \S_int[2] ;
 wire \S_int[3] ;
 wire \S_int[4] ;
 wire \S_int[5] ;
 wire \S_int[6] ;
 wire \S_int[7] ;
 wire \S_int[8] ;
 wire \S_int[9] ;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire clknet_0_CLK;
 wire clknet_2_0__leaf_CLK;
 wire clknet_2_1__leaf_CLK;
 wire clknet_2_2__leaf_CLK;
 wire clknet_2_3__leaf_CLK;

 sky130_fd_sc_hd__or2_1 _081_ (.A(\B_reg[15] ),
    .B(\A_reg[15] ),
    .X(_034_));
 sky130_fd_sc_hd__nor2_1 _082_ (.A(\B_reg[14] ),
    .B(\A_reg[14] ),
    .Y(_035_));
 sky130_fd_sc_hd__nor2_2 _083_ (.A(\B_reg[4] ),
    .B(\A_reg[4] ),
    .Y(_036_));
 sky130_fd_sc_hd__o22a_1 _084_ (.A1(\B_reg[7] ),
    .A2(\A_reg[7] ),
    .B1(\B_reg[6] ),
    .B2(\A_reg[6] ),
    .X(_037_));
 sky130_fd_sc_hd__or2_1 _085_ (.A(\B_reg[5] ),
    .B(\A_reg[5] ),
    .X(_038_));
 sky130_fd_sc_hd__nand2_1 _086_ (.A(_037_),
    .B(_038_),
    .Y(_039_));
 sky130_fd_sc_hd__nor2_1 _087_ (.A(\B_reg[3] ),
    .B(\A_reg[3] ),
    .Y(_040_));
 sky130_fd_sc_hd__nor2_1 _088_ (.A(\B_reg[2] ),
    .B(\A_reg[2] ),
    .Y(_041_));
 sky130_fd_sc_hd__or2_1 _089_ (.A(_040_),
    .B(_041_),
    .X(_042_));
 sky130_fd_sc_hd__or2_1 _090_ (.A(\B_reg[1] ),
    .B(\A_reg[1] ),
    .X(_043_));
 sky130_fd_sc_hd__a22o_1 _091_ (.A1(\B_reg[1] ),
    .A2(\A_reg[1] ),
    .B1(\B_reg[0] ),
    .B2(\A_reg[0] ),
    .X(_044_));
 sky130_fd_sc_hd__o221a_1 _092_ (.A1(\B_reg[1] ),
    .A2(\A_reg[1] ),
    .B1(\B_reg[0] ),
    .B2(\A_reg[0] ),
    .C1(CIN_reg),
    .X(_045_));
 sky130_fd_sc_hd__a21oi_1 _093_ (.A1(_043_),
    .A2(_044_),
    .B1(_045_),
    .Y(_046_));
 sky130_fd_sc_hd__nand2_1 _094_ (.A(\B_reg[2] ),
    .B(\A_reg[2] ),
    .Y(_047_));
 sky130_fd_sc_hd__nand2_1 _095_ (.A(\B_reg[3] ),
    .B(\A_reg[3] ),
    .Y(_048_));
 sky130_fd_sc_hd__o221a_2 _096_ (.A1(_042_),
    .A2(_046_),
    .B1(_047_),
    .B2(_040_),
    .C1(_048_),
    .X(_049_));
 sky130_fd_sc_hd__o211a_1 _097_ (.A1(\B_reg[7] ),
    .A2(\A_reg[7] ),
    .B1(\B_reg[6] ),
    .C1(\A_reg[6] ),
    .X(_050_));
 sky130_fd_sc_hd__a22o_1 _098_ (.A1(\B_reg[5] ),
    .A2(\A_reg[5] ),
    .B1(\B_reg[4] ),
    .B2(\A_reg[4] ),
    .X(_051_));
 sky130_fd_sc_hd__a32o_1 _099_ (.A1(_037_),
    .A2(_038_),
    .A3(_051_),
    .B1(\A_reg[7] ),
    .B2(\B_reg[7] ),
    .X(_052_));
 sky130_fd_sc_hd__nor2_1 _100_ (.A(_050_),
    .B(_052_),
    .Y(_053_));
 sky130_fd_sc_hd__o31ai_4 _101_ (.A1(_036_),
    .A2(_039_),
    .A3(_049_),
    .B1(_053_),
    .Y(_054_));
 sky130_fd_sc_hd__or2_1 _102_ (.A(\B_reg[8] ),
    .B(\A_reg[8] ),
    .X(_055_));
 sky130_fd_sc_hd__or2_1 _103_ (.A(\B_reg[10] ),
    .B(\A_reg[10] ),
    .X(_056_));
 sky130_fd_sc_hd__or2_1 _104_ (.A(\B_reg[11] ),
    .B(\A_reg[11] ),
    .X(_057_));
 sky130_fd_sc_hd__or2_1 _105_ (.A(\B_reg[9] ),
    .B(\A_reg[9] ),
    .X(_058_));
 sky130_fd_sc_hd__and3_1 _106_ (.A(_056_),
    .B(_057_),
    .C(_058_),
    .X(_059_));
 sky130_fd_sc_hd__nand2_1 _107_ (.A(\B_reg[9] ),
    .B(\A_reg[9] ),
    .Y(_060_));
 sky130_fd_sc_hd__nand2_1 _108_ (.A(\B_reg[8] ),
    .B(\A_reg[8] ),
    .Y(_061_));
 sky130_fd_sc_hd__nand2_1 _109_ (.A(_060_),
    .B(_061_),
    .Y(_062_));
 sky130_fd_sc_hd__nand2_1 _110_ (.A(\B_reg[10] ),
    .B(\A_reg[10] ),
    .Y(_063_));
 sky130_fd_sc_hd__a21bo_1 _111_ (.A1(_058_),
    .A2(_062_),
    .B1_N(_063_),
    .X(_064_));
 sky130_fd_sc_hd__and2_1 _112_ (.A(\B_reg[11] ),
    .B(\A_reg[11] ),
    .X(_065_));
 sky130_fd_sc_hd__a31o_1 _113_ (.A1(_056_),
    .A2(_057_),
    .A3(_064_),
    .B1(_065_),
    .X(_066_));
 sky130_fd_sc_hd__a31o_1 _114_ (.A1(_054_),
    .A2(_055_),
    .A3(_059_),
    .B1(_066_),
    .X(_067_));
 sky130_fd_sc_hd__or2_1 _115_ (.A(\B_reg[12] ),
    .B(\A_reg[12] ),
    .X(_068_));
 sky130_fd_sc_hd__o21a_1 _116_ (.A1(\B_reg[13] ),
    .A2(\A_reg[13] ),
    .B1(_068_),
    .X(_069_));
 sky130_fd_sc_hd__o211a_1 _117_ (.A1(\B_reg[13] ),
    .A2(\A_reg[13] ),
    .B1(\B_reg[12] ),
    .C1(\A_reg[12] ),
    .X(_070_));
 sky130_fd_sc_hd__a21o_1 _118_ (.A1(\B_reg[13] ),
    .A2(\A_reg[13] ),
    .B1(_070_),
    .X(_071_));
 sky130_fd_sc_hd__a21oi_1 _119_ (.A1(_067_),
    .A2(_069_),
    .B1(_071_),
    .Y(_072_));
 sky130_fd_sc_hd__nand2_1 _120_ (.A(\B_reg[14] ),
    .B(\A_reg[14] ),
    .Y(_073_));
 sky130_fd_sc_hd__o21ai_1 _121_ (.A1(_035_),
    .A2(_072_),
    .B1(_073_),
    .Y(_074_));
 sky130_fd_sc_hd__nand2_1 _122_ (.A(\B_reg[15] ),
    .B(\A_reg[15] ),
    .Y(_075_));
 sky130_fd_sc_hd__a21bo_1 _123_ (.A1(_034_),
    .A2(_074_),
    .B1_N(_075_),
    .X(\C[16] ));
 sky130_fd_sc_hd__o21ai_1 _124_ (.A1(\B_reg[0] ),
    .A2(\A_reg[0] ),
    .B1(CIN_reg),
    .Y(_076_));
 sky130_fd_sc_hd__nand2_1 _125_ (.A(\B_reg[0] ),
    .B(\A_reg[0] ),
    .Y(_077_));
 sky130_fd_sc_hd__or3_1 _126_ (.A(\B_reg[0] ),
    .B(\A_reg[0] ),
    .C(CIN_reg),
    .X(_078_));
 sky130_fd_sc_hd__and3_1 _127_ (.A(\B_reg[0] ),
    .B(\A_reg[0] ),
    .C(CIN_reg),
    .X(_079_));
 sky130_fd_sc_hd__a31o_1 _128_ (.A1(_076_),
    .A2(_077_),
    .A3(_078_),
    .B1(_079_),
    .X(\S_int[0] ));
 sky130_fd_sc_hd__nand2_1 _129_ (.A(_076_),
    .B(_077_),
    .Y(_080_));
 sky130_fd_sc_hd__nand2_1 _130_ (.A(\B_reg[1] ),
    .B(\A_reg[1] ),
    .Y(_000_));
 sky130_fd_sc_hd__and2_1 _131_ (.A(_043_),
    .B(_000_),
    .X(_001_));
 sky130_fd_sc_hd__xor2_1 _132_ (.A(_080_),
    .B(_001_),
    .X(\S_int[1] ));
 sky130_fd_sc_hd__and2b_1 _133_ (.A_N(_041_),
    .B(_047_),
    .X(_002_));
 sky130_fd_sc_hd__xnor2_1 _134_ (.A(_046_),
    .B(_002_),
    .Y(\S_int[2] ));
 sky130_fd_sc_hd__and2b_1 _135_ (.A_N(_040_),
    .B(_048_),
    .X(_003_));
 sky130_fd_sc_hd__nand2_1 _136_ (.A(_043_),
    .B(_044_),
    .Y(_004_));
 sky130_fd_sc_hd__or2b_1 _137_ (.A(_041_),
    .B_N(_045_),
    .X(_005_));
 sky130_fd_sc_hd__o211a_1 _138_ (.A1(_036_),
    .A2(_004_),
    .B1(_047_),
    .C1(_005_),
    .X(_006_));
 sky130_fd_sc_hd__xnor2_1 _139_ (.A(_003_),
    .B(_006_),
    .Y(\S_int[3] ));
 sky130_fd_sc_hd__and2_1 _140_ (.A(\B_reg[4] ),
    .B(\A_reg[4] ),
    .X(_007_));
 sky130_fd_sc_hd__nor2_1 _141_ (.A(_036_),
    .B(_007_),
    .Y(_008_));
 sky130_fd_sc_hd__xnor2_1 _142_ (.A(_049_),
    .B(_008_),
    .Y(\S_int[4] ));
 sky130_fd_sc_hd__nand2_1 _143_ (.A(\B_reg[5] ),
    .B(\A_reg[5] ),
    .Y(_009_));
 sky130_fd_sc_hd__nand2_1 _144_ (.A(_038_),
    .B(_009_),
    .Y(_010_));
 sky130_fd_sc_hd__nor2_1 _145_ (.A(_036_),
    .B(_049_),
    .Y(_011_));
 sky130_fd_sc_hd__or2_1 _146_ (.A(_007_),
    .B(_011_),
    .X(_012_));
 sky130_fd_sc_hd__xnor2_1 _147_ (.A(_010_),
    .B(_012_),
    .Y(\S_int[5] ));
 sky130_fd_sc_hd__nor2_1 _148_ (.A(\B_reg[6] ),
    .B(\A_reg[6] ),
    .Y(_013_));
 sky130_fd_sc_hd__nand2_1 _149_ (.A(\B_reg[6] ),
    .B(\A_reg[6] ),
    .Y(_014_));
 sky130_fd_sc_hd__and2b_1 _150_ (.A_N(_013_),
    .B(_014_),
    .X(_015_));
 sky130_fd_sc_hd__o21ai_1 _151_ (.A1(_051_),
    .A2(_011_),
    .B1(_038_),
    .Y(_016_));
 sky130_fd_sc_hd__xnor2_1 _152_ (.A(_015_),
    .B(_016_),
    .Y(\S_int[6] ));
 sky130_fd_sc_hd__xnor2_1 _153_ (.A(\B_reg[7] ),
    .B(\A_reg[7] ),
    .Y(_017_));
 sky130_fd_sc_hd__o21ai_1 _154_ (.A1(_013_),
    .A2(_016_),
    .B1(_014_),
    .Y(_018_));
 sky130_fd_sc_hd__xnor2_1 _155_ (.A(_017_),
    .B(_018_),
    .Y(\S_int[7] ));
 sky130_fd_sc_hd__nand2_1 _156_ (.A(_055_),
    .B(_061_),
    .Y(_019_));
 sky130_fd_sc_hd__xnor2_1 _157_ (.A(_054_),
    .B(_019_),
    .Y(\S_int[8] ));
 sky130_fd_sc_hd__nand2_1 _158_ (.A(_058_),
    .B(_060_),
    .Y(_020_));
 sky130_fd_sc_hd__a21bo_1 _159_ (.A1(_054_),
    .A2(_055_),
    .B1_N(_061_),
    .X(_021_));
 sky130_fd_sc_hd__xnor2_1 _160_ (.A(_020_),
    .B(_021_),
    .Y(\S_int[9] ));
 sky130_fd_sc_hd__nand2_1 _161_ (.A(_056_),
    .B(_063_),
    .Y(_022_));
 sky130_fd_sc_hd__a21o_1 _162_ (.A1(_054_),
    .A2(_055_),
    .B1(_062_),
    .X(_023_));
 sky130_fd_sc_hd__and2_1 _163_ (.A(_058_),
    .B(_023_),
    .X(_024_));
 sky130_fd_sc_hd__xnor2_1 _164_ (.A(_022_),
    .B(_024_),
    .Y(\S_int[10] ));
 sky130_fd_sc_hd__nand2_1 _165_ (.A(\B_reg[11] ),
    .B(\A_reg[11] ),
    .Y(_025_));
 sky130_fd_sc_hd__nand2_1 _166_ (.A(_057_),
    .B(_025_),
    .Y(_026_));
 sky130_fd_sc_hd__a21bo_1 _167_ (.A1(_056_),
    .A2(_024_),
    .B1_N(_063_),
    .X(_027_));
 sky130_fd_sc_hd__xnor2_1 _168_ (.A(_026_),
    .B(_027_),
    .Y(\S_int[11] ));
 sky130_fd_sc_hd__nand2_1 _169_ (.A(\B_reg[12] ),
    .B(\A_reg[12] ),
    .Y(_028_));
 sky130_fd_sc_hd__nand2_1 _170_ (.A(_068_),
    .B(_028_),
    .Y(_029_));
 sky130_fd_sc_hd__xnor2_1 _171_ (.A(_067_),
    .B(_029_),
    .Y(\S_int[12] ));
 sky130_fd_sc_hd__xnor2_1 _172_ (.A(\B_reg[13] ),
    .B(\A_reg[13] ),
    .Y(_030_));
 sky130_fd_sc_hd__a21bo_1 _173_ (.A1(_067_),
    .A2(_068_),
    .B1_N(_028_),
    .X(_031_));
 sky130_fd_sc_hd__xnor2_1 _174_ (.A(_030_),
    .B(_031_),
    .Y(\S_int[13] ));
 sky130_fd_sc_hd__and2b_1 _175_ (.A_N(_035_),
    .B(_073_),
    .X(_032_));
 sky130_fd_sc_hd__xnor2_1 _176_ (.A(_072_),
    .B(_032_),
    .Y(\S_int[14] ));
 sky130_fd_sc_hd__nand2_1 _177_ (.A(_034_),
    .B(_075_),
    .Y(_033_));
 sky130_fd_sc_hd__xnor2_1 _178_ (.A(_074_),
    .B(_033_),
    .Y(\S_int[15] ));
 sky130_fd_sc_hd__dfrtp_1 _179_ (.CLK(clknet_2_1__leaf_CLK),
    .D(\S_int[0] ),
    .RESET_B(net34),
    .Q(net36));
 sky130_fd_sc_hd__dfrtp_1 _180_ (.CLK(clknet_2_1__leaf_CLK),
    .D(\S_int[1] ),
    .RESET_B(net34),
    .Q(net43));
 sky130_fd_sc_hd__dfrtp_1 _181_ (.CLK(clknet_2_1__leaf_CLK),
    .D(\S_int[2] ),
    .RESET_B(net34),
    .Q(net44));
 sky130_fd_sc_hd__dfrtp_1 _182_ (.CLK(clknet_2_1__leaf_CLK),
    .D(\S_int[3] ),
    .RESET_B(net34),
    .Q(net45));
 sky130_fd_sc_hd__dfrtp_1 _183_ (.CLK(clknet_2_1__leaf_CLK),
    .D(\S_int[4] ),
    .RESET_B(net34),
    .Q(net46));
 sky130_fd_sc_hd__dfrtp_1 _184_ (.CLK(clknet_2_1__leaf_CLK),
    .D(\S_int[5] ),
    .RESET_B(net34),
    .Q(net47));
 sky130_fd_sc_hd__dfrtp_1 _185_ (.CLK(clknet_2_1__leaf_CLK),
    .D(\S_int[6] ),
    .RESET_B(net34),
    .Q(net48));
 sky130_fd_sc_hd__dfrtp_1 _186_ (.CLK(clknet_2_1__leaf_CLK),
    .D(\S_int[7] ),
    .RESET_B(net34),
    .Q(net49));
 sky130_fd_sc_hd__dfrtp_1 _187_ (.CLK(clknet_2_1__leaf_CLK),
    .D(\S_int[8] ),
    .RESET_B(net34),
    .Q(net50));
 sky130_fd_sc_hd__dfrtp_1 _188_ (.CLK(clknet_2_1__leaf_CLK),
    .D(\S_int[9] ),
    .RESET_B(net34),
    .Q(net51));
 sky130_fd_sc_hd__dfrtp_1 _189_ (.CLK(clknet_2_3__leaf_CLK),
    .D(\S_int[10] ),
    .RESET_B(net34),
    .Q(net37));
 sky130_fd_sc_hd__dfrtp_1 _190_ (.CLK(clknet_2_3__leaf_CLK),
    .D(\S_int[11] ),
    .RESET_B(net34),
    .Q(net38));
 sky130_fd_sc_hd__dfrtp_1 _191_ (.CLK(clknet_2_3__leaf_CLK),
    .D(\S_int[12] ),
    .RESET_B(net34),
    .Q(net39));
 sky130_fd_sc_hd__dfrtp_1 _192_ (.CLK(clknet_2_3__leaf_CLK),
    .D(\S_int[13] ),
    .RESET_B(net34),
    .Q(net40));
 sky130_fd_sc_hd__dfrtp_1 _193_ (.CLK(clknet_2_3__leaf_CLK),
    .D(\S_int[14] ),
    .RESET_B(net34),
    .Q(net41));
 sky130_fd_sc_hd__dfrtp_1 _194_ (.CLK(clknet_2_3__leaf_CLK),
    .D(\S_int[15] ),
    .RESET_B(net34),
    .Q(net42));
 sky130_fd_sc_hd__dfrtp_1 _195_ (.CLK(clknet_2_3__leaf_CLK),
    .D(\C[16] ),
    .RESET_B(net34),
    .Q(net35));
 sky130_fd_sc_hd__dfrtp_1 _196_ (.CLK(clknet_2_0__leaf_CLK),
    .D(net17),
    .RESET_B(net34),
    .Q(\B_reg[0] ));
 sky130_fd_sc_hd__dfrtp_1 _197_ (.CLK(clknet_2_0__leaf_CLK),
    .D(net24),
    .RESET_B(net34),
    .Q(\B_reg[1] ));
 sky130_fd_sc_hd__dfrtp_1 _198_ (.CLK(clknet_2_0__leaf_CLK),
    .D(net25),
    .RESET_B(net34),
    .Q(\B_reg[2] ));
 sky130_fd_sc_hd__dfrtp_1 _199_ (.CLK(clknet_2_0__leaf_CLK),
    .D(net26),
    .RESET_B(net34),
    .Q(\B_reg[3] ));
 sky130_fd_sc_hd__dfrtp_1 _200_ (.CLK(clknet_2_0__leaf_CLK),
    .D(net27),
    .RESET_B(net34),
    .Q(\B_reg[4] ));
 sky130_fd_sc_hd__dfrtp_1 _201_ (.CLK(clknet_2_0__leaf_CLK),
    .D(net28),
    .RESET_B(net34),
    .Q(\B_reg[5] ));
 sky130_fd_sc_hd__dfrtp_1 _202_ (.CLK(clknet_2_1__leaf_CLK),
    .D(net29),
    .RESET_B(net34),
    .Q(\B_reg[6] ));
 sky130_fd_sc_hd__dfrtp_1 _203_ (.CLK(clknet_2_1__leaf_CLK),
    .D(net30),
    .RESET_B(net34),
    .Q(\B_reg[7] ));
 sky130_fd_sc_hd__dfrtp_1 _204_ (.CLK(clknet_2_1__leaf_CLK),
    .D(net31),
    .RESET_B(net34),
    .Q(\B_reg[8] ));
 sky130_fd_sc_hd__dfrtp_1 _205_ (.CLK(clknet_2_1__leaf_CLK),
    .D(net32),
    .RESET_B(net34),
    .Q(\B_reg[9] ));
 sky130_fd_sc_hd__dfrtp_1 _206_ (.CLK(clknet_2_1__leaf_CLK),
    .D(net18),
    .RESET_B(net34),
    .Q(\B_reg[10] ));
 sky130_fd_sc_hd__dfrtp_1 _207_ (.CLK(clknet_2_1__leaf_CLK),
    .D(net19),
    .RESET_B(net34),
    .Q(\B_reg[11] ));
 sky130_fd_sc_hd__dfrtp_1 _208_ (.CLK(clknet_2_1__leaf_CLK),
    .D(net20),
    .RESET_B(net34),
    .Q(\B_reg[12] ));
 sky130_fd_sc_hd__dfrtp_1 _209_ (.CLK(clknet_2_3__leaf_CLK),
    .D(net21),
    .RESET_B(net34),
    .Q(\B_reg[13] ));
 sky130_fd_sc_hd__dfrtp_1 _210_ (.CLK(clknet_2_3__leaf_CLK),
    .D(net22),
    .RESET_B(net34),
    .Q(\B_reg[14] ));
 sky130_fd_sc_hd__dfrtp_1 _211_ (.CLK(clknet_2_3__leaf_CLK),
    .D(net23),
    .RESET_B(net34),
    .Q(\B_reg[15] ));
 sky130_fd_sc_hd__dfrtp_1 _212_ (.CLK(clknet_2_0__leaf_CLK),
    .D(net1),
    .RESET_B(net34),
    .Q(\A_reg[0] ));
 sky130_fd_sc_hd__dfrtp_1 _213_ (.CLK(clknet_2_0__leaf_CLK),
    .D(net8),
    .RESET_B(net34),
    .Q(\A_reg[1] ));
 sky130_fd_sc_hd__dfrtp_1 _214_ (.CLK(clknet_2_0__leaf_CLK),
    .D(net9),
    .RESET_B(net34),
    .Q(\A_reg[2] ));
 sky130_fd_sc_hd__dfrtp_1 _215_ (.CLK(clknet_2_0__leaf_CLK),
    .D(net10),
    .RESET_B(net34),
    .Q(\A_reg[3] ));
 sky130_fd_sc_hd__dfrtp_1 _216_ (.CLK(clknet_2_0__leaf_CLK),
    .D(net11),
    .RESET_B(net34),
    .Q(\A_reg[4] ));
 sky130_fd_sc_hd__dfrtp_1 _217_ (.CLK(clknet_2_0__leaf_CLK),
    .D(net12),
    .RESET_B(net34),
    .Q(\A_reg[5] ));
 sky130_fd_sc_hd__dfrtp_1 _218_ (.CLK(clknet_2_0__leaf_CLK),
    .D(net13),
    .RESET_B(net34),
    .Q(\A_reg[6] ));
 sky130_fd_sc_hd__dfrtp_1 _219_ (.CLK(clknet_2_2__leaf_CLK),
    .D(net14),
    .RESET_B(net34),
    .Q(\A_reg[7] ));
 sky130_fd_sc_hd__dfrtp_1 _220_ (.CLK(clknet_2_2__leaf_CLK),
    .D(net15),
    .RESET_B(net34),
    .Q(\A_reg[8] ));
 sky130_fd_sc_hd__dfrtp_1 _221_ (.CLK(clknet_2_2__leaf_CLK),
    .D(net16),
    .RESET_B(net34),
    .Q(\A_reg[9] ));
 sky130_fd_sc_hd__dfrtp_1 _222_ (.CLK(clknet_2_2__leaf_CLK),
    .D(net2),
    .RESET_B(net34),
    .Q(\A_reg[10] ));
 sky130_fd_sc_hd__dfrtp_1 _223_ (.CLK(clknet_2_2__leaf_CLK),
    .D(net3),
    .RESET_B(net34),
    .Q(\A_reg[11] ));
 sky130_fd_sc_hd__dfrtp_1 _224_ (.CLK(clknet_2_2__leaf_CLK),
    .D(net4),
    .RESET_B(net34),
    .Q(\A_reg[12] ));
 sky130_fd_sc_hd__dfrtp_1 _225_ (.CLK(clknet_2_2__leaf_CLK),
    .D(net5),
    .RESET_B(net34),
    .Q(\A_reg[13] ));
 sky130_fd_sc_hd__dfrtp_1 _226_ (.CLK(clknet_2_2__leaf_CLK),
    .D(net6),
    .RESET_B(net34),
    .Q(\A_reg[14] ));
 sky130_fd_sc_hd__dfrtp_1 _227_ (.CLK(clknet_2_2__leaf_CLK),
    .D(net7),
    .RESET_B(net34),
    .Q(\A_reg[15] ));
 sky130_fd_sc_hd__dfrtp_1 _228_ (.CLK(clknet_2_2__leaf_CLK),
    .D(net33),
    .RESET_B(net34),
    .Q(CIN_reg));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_116 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(A[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(A[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(A[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(A[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(A[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(A[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(A[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(A[1]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(A[2]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(A[3]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(A[4]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(A[5]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(A[6]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(A[7]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(A[8]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(A[9]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(B[0]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(B[10]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(B[11]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(B[12]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(B[13]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(B[14]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(B[15]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(B[1]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(B[2]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(B[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(B[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(B[5]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(B[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(B[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(B[8]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(B[9]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(CIN),
    .X(net33));
 sky130_fd_sc_hd__buf_12 input34 (.A(RST_N),
    .X(net34));
 sky130_fd_sc_hd__buf_1 output35 (.A(net35),
    .X(COUT));
 sky130_fd_sc_hd__clkbuf_1 output36 (.A(net36),
    .X(S[0]));
 sky130_fd_sc_hd__buf_1 output37 (.A(net37),
    .X(S[10]));
 sky130_fd_sc_hd__buf_1 output38 (.A(net38),
    .X(S[11]));
 sky130_fd_sc_hd__buf_1 output39 (.A(net39),
    .X(S[12]));
 sky130_fd_sc_hd__buf_1 output40 (.A(net40),
    .X(S[13]));
 sky130_fd_sc_hd__buf_1 output41 (.A(net41),
    .X(S[14]));
 sky130_fd_sc_hd__buf_1 output42 (.A(net42),
    .X(S[15]));
 sky130_fd_sc_hd__buf_1 output43 (.A(net43),
    .X(S[1]));
 sky130_fd_sc_hd__buf_1 output44 (.A(net44),
    .X(S[2]));
 sky130_fd_sc_hd__buf_1 output45 (.A(net45),
    .X(S[3]));
 sky130_fd_sc_hd__buf_1 output46 (.A(net46),
    .X(S[4]));
 sky130_fd_sc_hd__buf_1 output47 (.A(net47),
    .X(S[5]));
 sky130_fd_sc_hd__buf_1 output48 (.A(net48),
    .X(S[6]));
 sky130_fd_sc_hd__buf_1 output49 (.A(net49),
    .X(S[7]));
 sky130_fd_sc_hd__buf_1 output50 (.A(net50),
    .X(S[8]));
 sky130_fd_sc_hd__buf_1 output51 (.A(net51),
    .X(S[9]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_CLK (.A(CLK),
    .X(clknet_0_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_CLK (.A(clknet_0_CLK),
    .X(clknet_2_0__leaf_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_CLK (.A(clknet_0_CLK),
    .X(clknet_2_1__leaf_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_CLK (.A(clknet_0_CLK),
    .X(clknet_2_2__leaf_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_CLK (.A(clknet_0_CLK),
    .X(clknet_2_3__leaf_CLK));
 sky130_fd_sc_hd__bufinv_16 clkload0 (.A(clknet_2_0__leaf_CLK));
 sky130_fd_sc_hd__inv_6 clkload1 (.A(clknet_2_2__leaf_CLK));
 sky130_fd_sc_hd__inv_6 clkload2 (.A(clknet_2_3__leaf_CLK));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_141 ();
endmodule
